library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library lib;
use lib.textengine_package.all;

entity spriteengine_rom is
	port (clk : in std_logic);
end entity;

architecture x of spriteengine_rom is

begin

end architecture;
